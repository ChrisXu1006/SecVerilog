//=========================================================================
// Alternative Blocking Cache Control
//=========================================================================

`ifndef PLAB3_MEM_BLOCKING_CACHE_ALT_CTRL_V
`define PLAB3_MEM_BLOCKING_CACHE_ALT_CTRL_V

`include "plab5-mcore-define.v"
`include "plab3-mem-DecodeWben.v"
`include "vc-mem-msgs.v"
`include "vc-assert.v"

module plab3_mem_BlockingCacheAltCtrl
#(
  parameter size    = 256,            // Cache size in bytes

  parameter p_idx_shamt = 0,

  parameter p_opaque_nbits  = 8,

  // local parameters not meant to be set from outside
  parameter dbw     = 32,             // Short name for data bitwidth
  parameter abw     = 32,             // Short name for addr bitwidth
  parameter clw     = 128,            // Short name for cacheline bitwidth
  parameter nblocks = size*8/clw,     // Number of blocks in the cache

  parameter o = p_opaque_nbits
)
(
  input                                               clk,
  input                                               reset,

  // Cache Request

  inout												  cachereq_domain,
  input                                               cachereq_val,
  output reg                                          cachereq_rdy,

  // Cache Response

  output reg                                          cacheresp_val,
  input                                               cacheresp_rdy,

  // Memory Request

  output											  memreq_domain,
  output reg                                          memreq_val,
  input                                               memreq_rdy,

  // Memory Response

  input												  memresp_domain,
  input                                               memresp_val,
  output reg                                          memresp_rdy,

  // control signals (ctrl->dpath)
  output reg [1:0]                                    amo_sel,
  output reg                                          cachereq_en,
  output reg                                          memresp_en,
  output reg                                          is_refill,
  output reg                                          tag_array_0_wen,
  output reg                                          tag_array_0_ren,
  output reg                                          tag_array_1_wen,
  output reg                                          tag_array_1_ren,
  output                                              way_sel,
  output reg                                          data_array_wen,
  output reg                                          data_array_ren,
  // width of cacheline divided by number of bits per byte
  output reg [clw/8-1:0]                              data_array_wben,
  output reg                                          read_data_reg_en,
  output reg                                          read_tag_reg_en,
  output [$clog2(clw/dbw)-1:0]                        read_byte_sel,
  output reg [`VC_MEM_RESP_MSG_TYPE_NBITS(o,clw)-1:0] memreq_type,
  output reg [`VC_MEM_RESP_MSG_TYPE_NBITS(o,dbw)-1:0] cacheresp_type,

   // status signals (dpath->ctrl)
  input [`VC_MEM_REQ_MSG_TYPE_NBITS(o,abw,dbw)-1:0]   cachereq_type,
  input [`VC_MEM_REQ_MSG_ADDR_NBITS(o,abw,dbw)-1:0]   cachereq_addr,
  input                                               tag_match_0,
  input                                               tag_match_1,
  input												  nsbit_match_0,
  input												  nsbit_match_1
 );

  //----------------------------------------------------------------------
  // State Definitions
  //----------------------------------------------------------------------

  localparam STATE_IDLE						= 5'd0;
  localparam STATE_TAG_CHECK				= 5'd1;
  localparam STATE_READ_DATA_ACCESS			= 5'd2;
  localparam STATE_WRITE_DATA_ACCESS		= 5'd3;
  localparam STATE_WAIT						= 5'd4;
  localparam STATE_REFILL_REQUEST			= 5'd5;
  localparam STATE_REFILL_WAIT				= 5'd6;
  localparam STATE_REFILL_UPDATE			= 5'd7;
  localparam STATE_EVICT_PREPARE			= 5'd8;
  localparam STATE_EVICT_REQUEST			= 5'd9;
  localparam STATE_EVICT_WAIT				= 5'd10;
  localparam STATE_AMO_READ_DATA_ACCESS		= 5'd11;
  localparam STATE_AMO_WRITE_DATA_ACCESS	= 5'd12;
  localparam STATE_FAKE_READ_DATA_ACCESS	= 5'd13;
  localparam STATE_FAKE_WRITE_DATA_ACCESS	= 5'd14;
  localparam STATE_INIT_DATA_ACCESS			= 5'd15;

  //----------------------------------------------------------------------
  // State
  //----------------------------------------------------------------------

  always @( posedge clk ) begin
    if ( reset ) begin
      state_reg <= STATE_IDLE;
    end
    else begin
      state_reg <= state_next;
    end

	`ifdef DEBUG
		if ( state_reg === STATE_FAKE_READ_DATA_ACCESS )
			$display("enter fake read data access");
		else if ( state_reg === STATE_FAKE_WRITE_DATA_ACCESS )
			$display("enter fake write data access");
	`endif

  end

   //----------------------------------------------------------------------
  // State Transitions
  //----------------------------------------------------------------------

  wire in_go        = cachereq_val  && cachereq_rdy;
  wire out_go       = cacheresp_val && cacheresp_rdy;
  wire sec_0		= nsbit_match_0;
  wire sec_1		= nsbit_match_1;
  wire hit_0        = is_valid_0 && tag_match_0 && sec_0;
  wire hit_1        = is_valid_1 && tag_match_1 && sec_1;
  wire hit          = hit_0 || hit_1;
  wire fake_hit_0	= is_valid_0 && tag_match_0 && !sec_0;
  wire fake_hit_1	= is_valid_1 && tag_match_1 && !sec_1;
  wire fake_hit		= fake_hit_0 || fake_hit_1;
  wire is_read      = cachereq_type == `VC_MEM_REQ_MSG_TYPE_READ;
  wire is_write     = cachereq_type == `VC_MEM_REQ_MSG_TYPE_WRITE;
  wire is_init      = cachereq_type == `VC_MEM_REQ_MSG_TYPE_WRITE_INIT;
  wire is_amo       = amo_sel != 0;
  wire read_hit     = is_read && hit;
  wire fread_hit	= is_read && fake_hit;
  wire write_hit    = is_write && hit;
  wire fwrite_hit	= is_write && fake_hit;
  wire amo_hit      = is_amo && hit;
  wire miss_0       = !hit_0;
  wire miss_1       = !hit_1;
  wire refill       = (miss_0 && !is_dirty_0 && !lru_way) || (miss_1 && !is_dirty_1 && lru_way);
  wire evict        = (miss_0 && is_dirty_0 && !lru_way) || (miss_1 && is_dirty_1 && lru_way);

  reg [4:0] state_reg;
  reg [4:0] state_next;

  always @(*) begin

    state_next = state_reg;
    case ( state_reg )

      STATE_IDLE:
             if ( in_go        ) state_next = STATE_TAG_CHECK;

      STATE_TAG_CHECK:
             if ( is_init      ) state_next = STATE_INIT_DATA_ACCESS;
        else if ( read_hit     ) state_next = STATE_READ_DATA_ACCESS;
		else if ( fread_hit	   ) state_next = STATE_FAKE_READ_DATA_ACCESS;
        else if ( write_hit    ) state_next = STATE_WRITE_DATA_ACCESS;
		else if ( fwrite_hit   ) state_next = STATE_FAKE_WRITE_DATA_ACCESS;
        else if ( amo_hit      ) state_next = STATE_AMO_READ_DATA_ACCESS;
        else if ( refill       ) state_next = STATE_REFILL_REQUEST;
        else if ( evict        ) state_next = STATE_EVICT_PREPARE;

      STATE_READ_DATA_ACCESS:
        state_next = STATE_WAIT;

	  STATE_FAKE_READ_DATA_ACCESS:
		state_next = STATE_WAIT;

      STATE_WRITE_DATA_ACCESS:
        state_next = STATE_WAIT;

	  STATE_FAKE_WRITE_DATA_ACCESS:
		state_next = STATE_WAIT;

      STATE_INIT_DATA_ACCESS:
        state_next = STATE_WAIT;

      STATE_AMO_READ_DATA_ACCESS:
        state_next = STATE_AMO_WRITE_DATA_ACCESS;

      STATE_AMO_WRITE_DATA_ACCESS:
        state_next = STATE_WAIT;

      STATE_REFILL_REQUEST:
             if ( memreq_rdy   ) state_next = STATE_REFILL_WAIT;
        else if ( !memreq_rdy  ) state_next = STATE_REFILL_REQUEST;

      STATE_REFILL_WAIT:
             if ( memresp_val  ) state_next = STATE_REFILL_UPDATE;
        else if ( !memresp_val ) state_next = STATE_REFILL_WAIT;

      STATE_REFILL_UPDATE:
             if ( is_read  && memresp_domain <= cachereq_domain   ) 
								 state_next = STATE_READ_DATA_ACCESS;
		else if ( is_read  && memresp_domain >  cachereq_domain   )
								 state_next = STATE_FAKE_READ_DATA_ACCESS;
        else if ( is_write && memresp_domain <= cachereq_domain   ) 
								 state_next = STATE_WRITE_DATA_ACCESS;
		else if ( is_write && memresp_domain > cachereq_domain )
								 state_next = STATE_FAKE_WRITE_DATA_ACCESS;	
        else if ( is_amo       ) state_next = STATE_AMO_READ_DATA_ACCESS;

      STATE_EVICT_PREPARE:
        state_next = STATE_EVICT_REQUEST;

      STATE_EVICT_REQUEST:
             if ( memreq_rdy   ) state_next = STATE_EVICT_WAIT;
        else if ( !memreq_rdy  ) state_next = STATE_EVICT_REQUEST;

      STATE_EVICT_WAIT:
             if ( memresp_val  ) state_next = STATE_REFILL_REQUEST;
        else if ( !memresp_val ) state_next = STATE_EVICT_WAIT;

      STATE_WAIT:
             if ( out_go       ) state_next = STATE_IDLE;

    endcase

  end

  //----------------------------------------------------------------------
  // Valid/Dirty bits record
  //----------------------------------------------------------------------

  wire [2:0] cachereq_idx = cachereq_addr[4+p_idx_shamt +: 3];
  reg        valid_bit_in;
  reg        valid_bits_write_en;
  wire       valid_bits_write_en_0 = valid_bits_write_en && !way_sel;
  wire       valid_bits_write_en_1 = valid_bits_write_en && way_sel;
  wire       is_valid_0;
  wire       is_valid_1;

  vc_ResetRegfile_1r1w#(1,8) valid_bits_0
  (
    .clk        (clk),
    .reset      (reset),
    .read_addr  (cachereq_idx),
    .read_data  (is_valid_0),
    .write_en   (valid_bits_write_en_0),
    .write_addr (cachereq_idx),
    .write_data (valid_bit_in)
  );

  vc_ResetRegfile_1r1w#(1,8) valid_bits_1
  (
    .clk        (clk),
    .reset      (reset),
    .read_addr  (cachereq_idx),
    .read_data  (is_valid_1),
    .write_en   (valid_bits_write_en_1),
    .write_addr (cachereq_idx),
    .write_data (valid_bit_in)
  );

  reg        dirty_bit_in;
  reg        dirty_bits_write_en;
  wire       dirty_bits_write_en_0 = dirty_bits_write_en && !way_sel;
  wire       dirty_bits_write_en_1 = dirty_bits_write_en && way_sel;
  wire       is_dirty_0;
  wire       is_dirty_1;

  vc_ResetRegfile_1r1w#(1,8) dirty_bits_0
  (
    .clk        (clk),
    .reset      (reset),
    .read_addr  (cachereq_idx),
    .read_data  (is_dirty_0),
    .write_en   (dirty_bits_write_en_0),
    .write_addr (cachereq_idx),
    .write_data (dirty_bit_in)
  );

  vc_ResetRegfile_1r1w#(1,8) dirty_bits_1
  (
    .clk        (clk),
    .reset      (reset),
    .read_addr  (cachereq_idx),
    .read_data  (is_dirty_1),
    .write_en   (dirty_bits_write_en_1),
    .write_addr (cachereq_idx),
    .write_data (dirty_bit_in)
  );

  reg        lru_bit_in;
  reg        lru_bits_write_en;
  wire       lru_way;

  vc_ResetRegfile_1r1w#(1,8) lru_bits
  (
    .clk        (clk),
    .reset      (reset),
    .read_addr  (cachereq_idx),
    .read_data  (lru_way),
    .write_en   (lru_bits_write_en),
    .write_addr (cachereq_idx),
    .write_data (lru_bit_in)
  );

  //----------------------------------------------------------------------
  // Way selection.
  //   The way is determined in the tag check state, and is
  //   then recorded for the entire transaction
  //----------------------------------------------------------------------

  reg        way_record_en;
  reg        way_record_in;

  always @(*) begin
    if (hit) begin
      way_record_in = hit_0 ? 1'b0 :
                      ( hit_1 ? 1'b1 : 1'bx );
    end
    else
      way_record_in = lru_way; // If miss, write to the LRU way
  end

  vc_EnResetReg #(1, 0) way_record
  (
    .clk    (clk),
    .reset  (reset),
    .en     (way_record_en),
    .d      (way_record_in),
    .q      (way_sel)
  );

  //----------------------------------------------------------------------
  // State Outputs
  //----------------------------------------------------------------------

  reg tag_array_wen;
  reg tag_array_ren;

  always@(*) begin
	
	cachereq_rdy        = 1'b0;
	cacheresp_val       = 1'b0;
	memreq_val          = 1'b0;
    memresp_rdy         = 1'b0;
    cachereq_en         = 1'bx;
    memresp_en          = 1'bx;
    is_refill           = 1'bx;
    tag_array_wen       = 1'b0;
    tag_array_ren       = 1'b0;
	data_array_wen      = 1'b0;
    data_array_ren      = 1'b0;
    read_data_reg_en    = 1'b0;
    read_tag_reg_en     = 1'b0;
    memreq_type         = 1'bx;
    valid_bit_in        = 1'bx;
    valid_bits_write_en = 1'b0;
    dirty_bit_in        = 1'bx;
    dirty_bits_write_en = 1'b0;
    lru_bits_write_en   = 1'b0;
    way_record_en       = 1'b0;

	
	case ( state_reg )
		
		STATE_IDLE:	begin
			cachereq_rdy        = 1'b1;
			cacheresp_val       = 1'b0;
			memreq_val          = 1'b0;
    		memresp_rdy         = 1'b0;
    		cachereq_en         = 1'b1;
    		memresp_en          = 1'b0;
    		is_refill           = 1'bx;
    		tag_array_wen       = 1'b0;
    		tag_array_ren       = 1'b0;
    		data_array_wen      = 1'b0;
    		data_array_ren      = 1'b0;
    		read_data_reg_en    = 1'b0;
    		read_tag_reg_en     = 1'b0;
    		memreq_type         = 1'bx;
    		valid_bit_in        = 1'bx;
    		valid_bits_write_en = 1'b0;
    		dirty_bit_in        = 1'bx;
    		dirty_bits_write_en = 1'b0;
    		lru_bits_write_en   = 1'b0;
    		way_record_en       = 1'b0;
		end

		STATE_TAG_CHECK: begin
			cachereq_rdy        = 1'b0;
			cacheresp_val       = 1'b0;
			memreq_val          = 1'b0;
    		memresp_rdy         = 1'b0;
    		cachereq_en         = 1'b0;
    		memresp_en          = 1'b0;
    		is_refill           = 1'bx;
    		tag_array_wen       = 1'b0;
    		tag_array_ren       = 1'b1;
    		data_array_wen      = 1'b0;
    		data_array_ren      = 1'b0;
    		read_data_reg_en    = 1'b0;
    		read_tag_reg_en     = 1'b0;
    		memreq_type         = 1'bx;
    		valid_bit_in        = 1'bx;
    		valid_bits_write_en = 1'b0;
    		dirty_bit_in        = 1'bx;
    		dirty_bits_write_en = 1'b0;
    		lru_bits_write_en   = 1'b0;
    		way_record_en       = 1'b1;
		end

		STATE_READ_DATA_ACCESS: begin
			cachereq_rdy        = 1'b0;
			cacheresp_val       = 1'b0;
			memreq_val          = 1'b0;
    		memresp_rdy         = 1'b0;
    		cachereq_en         = 1'b0;
    		memresp_en          = 1'b0;
    		is_refill           = 1'bx;
    		tag_array_wen       = 1'b0;
    		tag_array_ren       = 1'b0;
    		data_array_wen      = 1'b0;
    		data_array_ren      = 1'b1;
    		read_data_reg_en    = 1'b1;
    		read_tag_reg_en     = 1'b0;
    		memreq_type         = 1'bx;
    		valid_bit_in        = 1'bx;
    		valid_bits_write_en = 1'b0;
    		dirty_bit_in        = 1'bx;
    		dirty_bits_write_en = 1'b0;
    		lru_bits_write_en   = 1'b1;
    		way_record_en       = 1'b0;
		end

		STATE_FAKE_READ_DATA_ACCESS: begin
			cachereq_rdy        = 1'b0;
			cacheresp_val       = 1'b0;
			memreq_val          = 1'b0;
    		memresp_rdy         = 1'b0;
    		cachereq_en         = 1'b0;
    		memresp_en          = 1'b0;
    		is_refill           = 1'bx;
    		tag_array_wen       = 1'b0;
    		tag_array_ren       = 1'b0;
    		data_array_wen      = 1'b0;
    		data_array_ren      = 1'b0;
    		read_data_reg_en    = 1'b1;
    		read_tag_reg_en     = 1'b0;
    		memreq_type         = 1'bx;
    		valid_bit_in        = 1'bx;
    		valid_bits_write_en = 1'b0;
    		dirty_bit_in        = 1'bx;
    		dirty_bits_write_en = 1'b0;
    		lru_bits_write_en   = 1'b0;
    		way_record_en       = 1'b0;
		end
		
		STATE_WRITE_DATA_ACCESS: begin
			cachereq_rdy        = 1'b0;
			cacheresp_val       = 1'b0;
			memreq_val          = 1'b0;
    		memresp_rdy         = 1'b0;
    		cachereq_en         = 1'b0;
    		memresp_en          = 1'b0;
    		is_refill           = 1'b0;
    		tag_array_wen       = 1'b1;
    		tag_array_ren       = 1'b0;
    		data_array_wen      = 1'b1;
    		data_array_ren      = 1'b0;
    		read_data_reg_en    = 1'b0;
    		read_tag_reg_en     = 1'b0;
    		memreq_type         = 1'bx;
    		valid_bit_in        = 1'b1;
    		valid_bits_write_en = 1'b1;
    		dirty_bit_in        = 1'b1;
    		dirty_bits_write_en = 1'b1;
    		lru_bits_write_en   = 1'b1;
    		way_record_en       = 1'b0;
		end

		STATE_FAKE_WRITE_DATA_ACCESS: begin
			cachereq_rdy        = 1'b0;
			cacheresp_val       = 1'b0;
			memreq_val          = 1'b0;
    		memresp_rdy         = 1'b0;
    		cachereq_en         = 1'b0;
    		memresp_en          = 1'b0;
    		is_refill           = 1'b0;
    		tag_array_wen       = 1'b0;
    		tag_array_ren       = 1'b0;
    		data_array_wen      = 1'b0;
    		data_array_ren      = 1'b0;
    		read_data_reg_en    = 1'b0;
    		read_tag_reg_en     = 1'b0;
    		memreq_type         = 1'bx;
    		valid_bit_in        = 1'bx;
    		valid_bits_write_en = 1'b0;
    		dirty_bit_in        = 1'bx;
    		dirty_bits_write_en = 1'b0;
    		lru_bits_write_en   = 1'b0;
    		way_record_en       = 1'b0;
		end

		STATE_INIT_DATA_ACCESS: begin
			cachereq_rdy        = 1'b0;
			cacheresp_val       = 1'b0;
			memreq_val          = 1'b0;
    		memresp_rdy         = 1'b0;
    		cachereq_en         = 1'b0;
    		memresp_en          = 1'b0;
    		is_refill           = 1'b0;
    		tag_array_wen       = 1'b1;
    		tag_array_ren       = 1'b0;
    		data_array_wen      = 1'b1;
    		data_array_ren      = 1'b0;
    		read_data_reg_en    = 1'b0;
    		read_tag_reg_en     = 1'b0;
    		memreq_type         = 1'bx;
    		valid_bit_in        = 1'b1;
    		valid_bits_write_en = 1'b1;
    		dirty_bit_in        = 1'b0;
    		dirty_bits_write_en = 1'b1;
    		lru_bits_write_en   = 1'b1;
    		way_record_en       = 1'b0;
		end

		STATE_AMO_READ_DATA_ACCESS: begin
			cachereq_rdy        = 1'b0;
			cacheresp_val       = 1'b0;
			memreq_val          = 1'b0;
    		memresp_rdy         = 1'b0;
    		cachereq_en         = 1'b0;
    		memresp_en          = 1'b0;
    		is_refill           = 1'bx;
    		tag_array_wen       = 1'b0;
    		tag_array_ren       = 1'b0;
    		data_array_wen      = 1'b0;
    		data_array_ren      = 1'b1;
    		read_data_reg_en    = 1'b1;
    		read_tag_reg_en     = 1'b0;
    		memreq_type         = 1'bx;
    		valid_bit_in        = 1'bx;
    		valid_bits_write_en = 1'b0;
    		dirty_bit_in        = 1'bx;
    		dirty_bits_write_en = 1'b0;
    		lru_bits_write_en   = 1'b1;
    		way_record_en       = 1'b0;
		end

		STATE_AMO_WRITE_DATA_ACCESS: begin
			cachereq_rdy        = 1'b0;
			cacheresp_val       = 1'b0;
			memreq_val          = 1'b0;
    		memresp_rdy         = 1'b0;
    		cachereq_en         = 1'b0;
    		memresp_en          = 1'b0;
    		is_refill           = 1'b0;
    		tag_array_wen       = 1'b1;
    		tag_array_ren       = 1'b0;
    		data_array_wen      = 1'b1;
    		data_array_ren      = 1'b0;
    		read_data_reg_en    = 1'b0;
    		read_tag_reg_en     = 1'b0;
    		memreq_type         = 1'bx;
    		valid_bit_in        = 1'b1;
    		valid_bits_write_en = 1'b1;
    		dirty_bit_in        = 1'b1;
    		dirty_bits_write_en = 1'b1;
    		lru_bits_write_en   = 1'b1;
    		way_record_en       = 1'b0;
		end

		STATE_REFILL_REQUEST: begin
			cachereq_rdy        = 1'b0;
			cacheresp_val       = 1'b0;
			memreq_val          = 1'b1;
    		memresp_rdy         = 1'b0;
    		cachereq_en         = 1'b0;
    		memresp_en          = 1'b0;
    		is_refill           = 1'bx;
    		tag_array_wen       = 1'b0;
    		tag_array_ren       = 1'b0;
    		data_array_wen      = 1'b0;
    		data_array_ren      = 1'b0;
    		read_data_reg_en    = 1'b0;
    		read_tag_reg_en     = 1'b0;
    		memreq_type         = 1'b0;
    		valid_bit_in        = 1'bx;
    		valid_bits_write_en = 1'b0;
    		dirty_bit_in        = 1'bx;
    		dirty_bits_write_en = 1'b0;
    		lru_bits_write_en   = 1'b0;
    		way_record_en       = 1'b0;
		end

		STATE_REFILL_WAIT: begin
			cachereq_rdy        = 1'b0;
			cacheresp_val       = 1'b0;
			memreq_val          = 1'b0;
    		memresp_rdy         = 1'b1;
    		cachereq_en         = 1'b0;
    		memresp_en          = 1'b1;
    		is_refill           = 1'bx;
    		tag_array_wen       = 1'b0;
    		tag_array_ren       = 1'b0;
    		data_array_wen      = 1'b0;
    		data_array_ren      = 1'b0;
    		read_data_reg_en    = 1'b0;
    		read_tag_reg_en     = 1'b0;
    		memreq_type         = 1'bx;
    		valid_bit_in        = 1'bx;
    		valid_bits_write_en = 1'b0;
    		dirty_bit_in        = 1'bx;
    		dirty_bits_write_en = 1'b0;
    		lru_bits_write_en   = 1'b0;
    		way_record_en       = 1'b0;
		end

		STATE_REFILL_UPDATE: begin
			cachereq_rdy        = 1'b0;
			cacheresp_val       = 1'b0;
			memreq_val          = 1'b0;
    		memresp_rdy         = 1'b0;
    		cachereq_en         = 1'b0;
    		memresp_en          = 1'b0;
    		is_refill           = 1'b1;
    		tag_array_wen       = 1'b1;
    		tag_array_ren       = 1'b0;
    		data_array_wen      = 1'b1;
    		data_array_ren      = 1'b0;
    		read_data_reg_en    = 1'b0;
    		read_tag_reg_en     = 1'b0;
    		memreq_type         = 1'bx;
    		valid_bit_in        = 1'b1;
    		valid_bits_write_en = 1'b1;
    		dirty_bit_in        = 1'b0;
    		dirty_bits_write_en = 1'b1;
    		lru_bits_write_en   = 1'b0;
    		way_record_en       = 1'b0;
		end

		STATE_EVICT_PREPARE: begin
			cachereq_rdy        = 1'b0;
			cacheresp_val       = 1'b0;
			memreq_val          = 1'b0;
    		memresp_rdy         = 1'b0;
    		cachereq_en         = 1'b0;
    		memresp_en          = 1'b0;
    		is_refill           = 1'bx;
    		tag_array_wen       = 1'b0;
    		tag_array_ren       = 1'b1;
    		data_array_wen      = 1'b0;
    		data_array_ren      = 1'b1;
    		read_data_reg_en    = 1'b1;
    		read_tag_reg_en     = 1'b1;
    		memreq_type         = 1'bx;
    		valid_bit_in        = 1'bx;
    		valid_bits_write_en = 1'b0;
    		dirty_bit_in        = 1'bx;
    		dirty_bits_write_en = 1'b0;
    		lru_bits_write_en   = 1'b0;
    		way_record_en       = 1'b0;
		end

		STATE_EVICT_REQUEST: begin
			cachereq_rdy        = 1'b0;
			cacheresp_val       = 1'b0;
			memreq_val          = 1'b1;
    		memresp_rdy         = 1'b0;
    		cachereq_en         = 1'b0;
    		memresp_en          = 1'b0;
    		is_refill           = 1'bx;
    		tag_array_wen       = 1'b0;
    		tag_array_ren       = 1'b0;
    		data_array_wen      = 1'b0;
    		data_array_ren      = 1'b0;
    		read_data_reg_en    = 1'b0;
    		read_tag_reg_en     = 1'b0;
    		memreq_type         = 1'b1;
    		valid_bit_in        = 1'bx;
    		valid_bits_write_en = 1'b0;
    		dirty_bit_in        = 1'bx;
    		dirty_bits_write_en = 1'b0;
    		lru_bits_write_en   = 1'b0;
    		way_record_en       = 1'b0;
		end

		STATE_EVICT_WAIT: begin
			cachereq_rdy        = 1'b0;
			cacheresp_val       = 1'b0;
			memreq_val          = 1'b0;
    		memresp_rdy         = 1'b1;
    		cachereq_en         = 1'b0;
    		memresp_en          = 1'b0;
    		is_refill           = 1'bx;
    		tag_array_wen       = 1'b0;
    		tag_array_ren       = 1'b0;
    		data_array_wen      = 1'b0;
    		data_array_ren      = 1'b0;
    		read_data_reg_en    = 1'b0;
    		read_tag_reg_en     = 1'b0;
    		memreq_type         = 1'bx;
    		valid_bit_in        = 1'bx;
    		valid_bits_write_en = 1'b0;
    		dirty_bit_in        = 1'bx;
    		dirty_bits_write_en = 1'b0;
    		lru_bits_write_en   = 1'b0;
    		way_record_en       = 1'b0;
		end

		STATE_WAIT: begin
			cachereq_rdy        = 1'b0;
			cacheresp_val       = 1'b1;
			memreq_val          = 1'b0;
    		memresp_rdy         = 1'b1;
    		cachereq_en         = 1'b0;
    		memresp_en          = 1'b0;
    		is_refill           = 1'bx;
    		tag_array_wen       = 1'b0;
    		tag_array_ren       = 1'b0;
    		data_array_wen      = 1'b0;
    		data_array_ren      = 1'b0;
    		read_data_reg_en    = 1'b0;
    		read_tag_reg_en     = 1'b0;
    		memreq_type         = 1'bx;
    		valid_bit_in        = 1'bx;
    		valid_bits_write_en = 1'b0;
    		dirty_bit_in        = 1'bx;
    		dirty_bits_write_en = 1'b0;
    		lru_bits_write_en   = 1'b0;
    		way_record_en       = 1'b0;
		end
	endcase
  end

  // lru bit determination
  always @(*) begin
    lru_bit_in = !way_sel;
  end

  // tag array enables

  always @(*) begin
    tag_array_0_wen = tag_array_wen && !way_sel;
    tag_array_0_ren = tag_array_ren;
    tag_array_1_wen = tag_array_wen && way_sel;
    tag_array_1_ren = tag_array_ren;
  end

  // Building data_array_wben
  // This is in control because we want to facilitate more complex patterns
  //   when we want to start supporting subword accesses

  wire [1:0] cachereq_offset = cachereq_addr[3:2];
  wire [15:0] wben_decoder_out;

  plab3_mem_DecoderWben#(2) wben_decoder
  (
    .in  (cachereq_offset),
    .out (wben_decoder_out)
  );

  // Choose byte to read from cacheline based on what the offset was

  assign read_byte_sel = cachereq_offset;

  // Pass cache request domain to memory request domain
  assign memreq_domain = cachereq_domain;

  // determine amo type

  always @(*) begin
    case ( cachereq_type )
      `VC_MEM_REQ_MSG_TYPE_AMO_ADD: amo_sel = 2'h1;
      `VC_MEM_REQ_MSG_TYPE_AMO_AND: amo_sel = 2'h2;
      `VC_MEM_REQ_MSG_TYPE_AMO_OR : amo_sel = 2'h3;
      default                     : amo_sel = 2'h0;
    endcase
  end

  // managing the wben

  always @(*) begin
    // Logic to enable writing of the entire cacheline in case of refill and just one word for writes and init

    if ( is_refill )
      data_array_wben = 16'hffff;
    else
      data_array_wben = wben_decoder_out;

    // Managing the cache response type based on cache request type

    cacheresp_type = cachereq_type;
  end

  //----------------------------------------------------------------------
  // Assertions
  //----------------------------------------------------------------------

  always @( posedge clk ) begin
    if ( !reset ) begin
      `VC_ASSERT_NOT_X( cachereq_val  );
      `VC_ASSERT_NOT_X( cacheresp_rdy );
      `VC_ASSERT_NOT_X( memreq_rdy    );
      `VC_ASSERT_NOT_X( memresp_val   );
    end
  end

endmodule

`endif
